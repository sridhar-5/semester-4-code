module xorgate(
    input a,
    input b,
    output y
);

xor x1(y,a,b);
endmodule
